*Simulation Title
************************************************

*In hSpICe, nO cASe-seNsiTivE.

*Understand this file with other's file.

*MAY THE FORCE BE WITH YOUR CIRCUIT

********************Options**********************
*https://www.cnblogs.com/qiushuixiaozhanshi/p/6273206.html

****general
.OPTION	INGOLD=2
.OPTION	PARHIER=LOCAL
.option BRIEF = 0



****for spice
*.OPTION	ARTIST=2
*.OPTION	PSF=2
*.OPTION	RUNLVL=5
*.OPTION	ACCURATE=1
*.OPTION	REDEFSUB=1
*.OPTION	LIS_NEW=1
*.option    NOMOD = 1



********************Model*************************
*.LIB '<filepath> filename' entryname
.lib '/dir/model.sp' tt
.temp 25

*******************Parameter**********************
.param vvdd=1.1


*******************Force Global Power********************
*Find them in your prenetlist file, they should be at the beginning.
.GLOBAL VDD! Vpower!


VG00 VDD!       0   vvdd $ This line means VDD! is vvdd(1.1V) higher than 0(GND/GND!/GROUND).
*If Vpower! is generated by some circuit, so no need to provide.

********************Netlist*************************
.inc 'netlist.sp'

********************Force Input***************************
V000    Vac               0    1
V001    Vpwl              0    pwl t1 v1, t2 v2 
V002

*********************************************
C1145141919810 VDD! NET_1145141919810 5n    $ This line means VDD! and NET_1145141919810 are connected with a 5nF capacitor.
R1145141919810 0    NET_1145141919810 4

*********************Measure*****************
.tran 1000n 100u 

.op
.probe V(*)
.probe V(*) I(*)
.probe V(*) I(*) isub(*)







.end
