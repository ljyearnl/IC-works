*Simulation Title
************************************************

*In hSpICe, nO cASe-seNsiTivE.

*Understand this file with other's file.

*MAY THE FORCE BE WITH YOUR CIRCUIT

********************Options**********************


****general
.OPTION	INGOLD=2
.OPTION	PARHIER=LOCAL
.option BRIEF = 0
.OPTION MEASFILE=1
.OPTION MEASFAIL=1


****for spice
*.OPTION	ARTIST=2
*.OPTION	PSF=2
*.OPTION	RUNLVL=5
*.OPTION	ACCURATE=1
*.OPTION	REDEFSUB=1
*.OPTION	LIS_NEW=1
*.option    NOMOD = 1



********************Model*************************
*.LIB '<filepath> filename' entryname
.lib '/dir/model.sp' tt
.temp 25

*******************Parameter**********************
.param vvdd=1.1


*******************Force Global Power********************
*Find them in your prenetlist file, they should be at the beginning.
.GLOBAL VDD! Vpower!


VG00 VDD!       0   vvdd $ This line means VDD! is vvdd(1.1V) higher than 0(GND/GND!/GROUND).
*If Vpower! is generated by some circuit, so no need to provide.

********************Netlist*************************
.inc 'netlist.sp'

********************Force Input***************************
V000    Vac               0    1
V001    Vpwl              0    pwl t1 v1, t2 v2 
V002

*********************************************
C1145141919810 VDD! NET_1145141919810 5n    $ This line means VDD! and NET_1145141919810 are connected with a 5nF capacitor.
R1145141919810 0    NET_1145141919810 4

*********************Measure*****************
.tran 1000n 100u sweep data=var

.data var T2 T1 T0
+0 0 0
+0 0 1
+0 1 0
+0 1 1
+1 0 0
+1 0 1
+1 1 0
+1 1 1


.op
.probe V(*)
.probe V(*) I(*)
.probe V(*) I(*) isub(*)


.meas tran Tfall WHEN v(OUT) VAL='vvdd*0.5' fall=10

.meas tran Tper1 trig v(OUT) VAL='vvdd*0.5' td='Tfall+1n' rise=1 targ v(OSCOUT)  VAL='vvdd*0.5' td='Tfall+1n' rise=2

.meas tran Tpw1 trig v(OUT) VAL='vvdd*0.5' td='Tfall+1n' rise=1 targ v(OSCOUT)  VAL='vvdd*0.5' td='Tfall+1n' fall=1







*test phase margin and gain of AMP, only works in hspice simulator

V_AC  STB1  STB2 0 
.LSTB mode=single vsource=V_AC
.ac DEC 100 1 1G 

.probe V(*) I(*) isub(*) 
.probe ac LSTB(DB:lvf) LSTB(P:lvf)

.meas ac PM find LSTB(P) when LSTB(DB)=0
.meas ac GAIN max LSTB(DB)



.end
